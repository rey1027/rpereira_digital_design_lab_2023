module lrl_logic_bit(input logic a,b, output logic out);

	assign out = a>>b;
endmodule