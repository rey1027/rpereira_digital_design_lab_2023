module main_tb;
    
    reg A, B, C, D;
    wire [6:0] seg;
    
	 main dut(.A(A), .B(B), .C(C), .D(D), .seg(seg));
    
    
    reg clk = 0;
    always #10 clk = ~clk;
    
    
    initial begin
	 
    A = 0; B = 0; C = 0; D = 0;
    #20;
    A = 0; B = 0; C = 0; D = 1;
    #20;
    A = 0; B = 0; C = 1; D = 0;
    #20;
    A = 0; B = 0; C = 1; D = 1;
    #20;
    A = 0; B = 1; C = 0; D = 0;
    #20;
    A = 0; B = 1; C = 0; D = 1;
    #20;
    A = 0; B = 1; C = 1; D = 0;
    #20;
    A = 0; B = 1; C = 1; D = 1;
    #20;
    A = 1; B = 0; C = 0; D = 0;
    #20;
    A = 1; B = 0; C = 0; D = 1;
    #20;
    A = 1; B = 0; C = 1; D = 0;
    #20
    A = 1; B = 0; C = 1; D = 1;
    #20;
    A = 1; B = 1; C = 0; D = 0;
    #20;
    A = 1; B = 1; C = 0; D = 1;
    #20;
    A = 1; B = 1; C = 1; D = 0;
    #20;
    A = 1; B = 1; C = 1; D = 1;
    #20; $finish;
    end
    
    // Monitor
    always @(posedge clk) begin
        $display("Input: A=%b, B=%b, C=%b, D=%b, Output: seg=%b", A, B, C, D, seg);
    end
endmodule