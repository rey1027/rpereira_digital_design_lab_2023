module lrl_arithmetic_bit(input logic a,b, output logic out);

	assign out = a>>>b;
endmodule