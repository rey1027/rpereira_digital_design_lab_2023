module main_tb;

//logic [3:0] dir;
//logic [15:0] score = 0;
//logic [15:0] inmatrix[0:3][0:3];
//logic win;
//logic lose;
//logic clk;
//logic reset;
//logic move_up;
//logic move_down;
//logic move_left;
//logic move_right;

logic ar;
logic ab;
logic iz;
logic de;
logic clk;
logic rst;
logic win;
logic loss;
logic [15:0] outmatrix[3:0][3:0];
logic [6:0] s0;
logic [6:0] s1;
logic [6:0] s2;
logic [6:0] s3;
logic vgaclk;
logic hsync; 
logic vsync;
logic sync_b;
logic blank_b;
logic [7:0] r;
logic [7:0] g;
logic [7:0] b;


//game2048 fsm(clk,reset,move_up,move_down,move_left,move_right,dir);

//controller_game game(dir,score,inmatrix,score,win,lose,inmatrix);

main game(ar,ab,iz,de,clk,rst,win,loss,s0,s1,s2,s3,vgaclk,hsync,vsync,sync_b,blank_b,r,g,b);

initial begin

// Reset a estado inicial
rst = 1; #50
clk = 0; rst = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;

ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
clk = 0; ar = 0; #50;
de = 1; clk = 1; #50;
clk = 0; de = 0; #50;
iz = 1; clk = 1; #50;
iz = 0; clk = 0; #50;
ab = 1; clk = 1; #50;
ab = 0; clk = 0; #50;
ar = 1; clk = 1; #50;
rst = 1; #50;
clk = 0; ar = 0; #50;
end 

endmodule